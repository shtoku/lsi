`include "consts_train.vh"

module dense_inner_10 #(
    parameter integer DATA_WIDTH1 = `N_LEN,
    parameter integer DATA_WIDTH2 = `N_LEN,
    parameter integer OUT_WIDTH     = `N_LEN
  ) (
    input  wire clk,
    input  wire rst_n,
    input  wire [10*DATA_WIDTH1-1:0] d1,
    input  wire [10*DATA_WIDTH2-1:0] d2,
    output reg  [OUT_WIDTH-1:0] q
  );


  // ----------------------------------------
  genvar i;

  // reg result
  reg  [OUT_WIDTH-1:0] mul  [0:9];
  reg  [OUT_WIDTH-1:0] add1 [0:3];
  reg  [OUT_WIDTH-1:0] add2 [0:1];


  // ----------------------------------------
  // function fixed_multiply
  function [OUT_WIDTH-1:0] fixed_mul;
    input signed [DATA_WIDTH1-1:0] num1;
    input signed [DATA_WIDTH2-1:0] num2;

    reg [2*OUT_WIDTH-1:0] mul;
    begin
      mul = num1 * num2;
      fixed_mul = mul[`F_LEN +: OUT_WIDTH]; 
    end
  endfunction  


  // ----------------------------------------
  // fixed multiply
  generate
    for (i = 0; i < 10; i = i + 1) begin
      always @(posedge clk, negedge rst_n) begin
        if (~rst_n)
          mul[i] <= 0;
        else
          mul[i] <= fixed_mul(d1[i*DATA_WIDTH1 +: DATA_WIDTH1], d2[i*DATA_WIDTH2 +: DATA_WIDTH2]);
      end
    end
  endgenerate

  // first add
  always @(posedge clk, negedge rst_n) begin
    if (~rst_n) begin
      add1[0] <= 0;
      add1[1] <= 0;
      add1[2] <= 0;
    end else begin
      add1[0] <= mul[0] + mul[1] + mul[2];
      add1[1] <= mul[3] + mul[4] + mul[5];
      add1[2] <= mul[6] + mul[7] + mul[8];
      add1[3] <= mul[9];
    end
  end

  // second add
  always @(posedge clk, negedge rst_n) begin
    if (~rst_n) begin
      add2[0] <= 0;
      add2[1] <= 0;
    end else begin
      add2[0] <= add1[0] + add1[1];
      add2[1] <= add1[2] + add1[3];
    end
  end

  // ouput add
  always @(posedge clk, negedge rst_n) begin
    if (~rst_n) begin
      q <= 0;
    end else begin
      q <= add2[0] + add2[1];
    end
  end
  
endmodule