`include "consts.vh"

module inner_24_tb ();

  reg clk;
  reg rst_n;
  reg run;
  reg signed [24*`N_LEN - 1:0] d1;
  reg signed [24*`N_LEN - 1:0] d2;
  wire signed [`N_LEN - 1:0] q;

  inner_24 inner_24_inst(clk, rst_n, run, d1, d2, q);

  initial clk = 0;
  always #5 clk = ~clk;

  initial begin
    $dumpvars;
    rst_n=0; run=0; //d1={{12{6'd1, 10'd0}}, {12{6'd1, 10'd0}}}; d2={{12{6'd1, 10'd0}}, {12{6'd1, 10'd0}}}; #10
    d1 = {
        16'b1111100111001110,
        16'b1111110010100101,
        16'b1111100100101111,
        16'b1111100010111110,
        16'b0000010111010110,
        16'b0000011101100010,
        16'b0000000100100000,
        16'b0000000010010110,
        16'b0000010000010110,
        16'b1111100010100111,
        16'b0000001110101011,
        16'b0000010011101111,
        16'b0000001000100011,
        16'b1111111000010100,
        16'b1111100101001000,
        16'b0000011100110110,
        16'b1111101011111100,
        16'b1111111000100110,
        16'b1111101101111000,
        16'b1111111011101001,
        16'b0000001000110111,
        16'b0000001010100101,
        16'b1111110101101011,
        16'b1111110000110101
    };
    d2 = {
        16'b0000000100011111,
        16'b1111111101010011,
        16'b0000001000000111,
        16'b1111110100101011,
        16'b0000001001011101,
        16'b1111111010100110,
        16'b0000000110001110,
        16'b1111111100001010,
        16'b1111111000110110,
        16'b0000001011110110,
        16'b1111111010001011,
        16'b1111111001111001,
        16'b1111111001111100,
        16'b0000000100011100,
        16'b1111111001111110,
        16'b0000001101000000,
        16'b0000000100010100,
        16'b0000000111000001,
        16'b1111111001001011,
        16'b0000000110000101,
        16'b1111111110111110,
        16'b1111111001000000,
        16'b1111110110011011,
        16'b0000000111111000
    }; #10
    rst_n=1; #10
    run=1; #10
    #300
    $finish;
  end

endmodule


//  1.5  => {6'b0000_01, 10'b10_0000_0000}
// -1.5  => {6'b1111_10, 10'b10_0000_0000}
// -1.25 => {6'b1111_10, 10'b11_0000_0000}